module myModule();
    initial
    begin
    $display("Hello World!"); // This will display a message
    $finish ; // This causes the simulation to end. Without, it would go on..and on.
    end
endmodule